// Verilog netlist created by TD v4.5.12562
// Sat Apr  4 21:26:26 2020

`timescale 1ns / 1ps
module mem  // al_ip/mem.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [16:0] addra;  // al_ip/mem.v(18)
  input clka;  // al_ip/mem.v(19)
  input rsta;  // al_ip/mem.v(20)
  output [7:0] doa;  // al_ip/mem.v(16)

  wire [0:3] addra_piped;
  wire  \inst_doa_mux_b0/B0_0 ;
  wire  \inst_doa_mux_b0/B0_1 ;
  wire  \inst_doa_mux_b0/B0_2 ;
  wire  \inst_doa_mux_b0/B0_3 ;
  wire  \inst_doa_mux_b0/B0_4 ;
  wire  \inst_doa_mux_b0/B0_5 ;
  wire  \inst_doa_mux_b0/B0_6 ;
  wire  \inst_doa_mux_b0/B0_7 ;
  wire  \inst_doa_mux_b0/B1_0 ;
  wire  \inst_doa_mux_b0/B1_1 ;
  wire  \inst_doa_mux_b0/B1_2 ;
  wire  \inst_doa_mux_b0/B1_3 ;
  wire  \inst_doa_mux_b0/B2_0 ;
  wire  \inst_doa_mux_b0/B2_1 ;
  wire  \inst_doa_mux_b1/B0_0 ;
  wire  \inst_doa_mux_b1/B0_1 ;
  wire  \inst_doa_mux_b1/B0_2 ;
  wire  \inst_doa_mux_b1/B0_3 ;
  wire  \inst_doa_mux_b1/B0_4 ;
  wire  \inst_doa_mux_b1/B0_5 ;
  wire  \inst_doa_mux_b1/B0_6 ;
  wire  \inst_doa_mux_b1/B0_7 ;
  wire  \inst_doa_mux_b1/B1_0 ;
  wire  \inst_doa_mux_b1/B1_1 ;
  wire  \inst_doa_mux_b1/B1_2 ;
  wire  \inst_doa_mux_b1/B1_3 ;
  wire  \inst_doa_mux_b1/B2_0 ;
  wire  \inst_doa_mux_b1/B2_1 ;
  wire  \inst_doa_mux_b2/B0_0 ;
  wire  \inst_doa_mux_b2/B0_1 ;
  wire  \inst_doa_mux_b2/B0_2 ;
  wire  \inst_doa_mux_b2/B0_3 ;
  wire  \inst_doa_mux_b2/B0_4 ;
  wire  \inst_doa_mux_b2/B0_5 ;
  wire  \inst_doa_mux_b2/B0_6 ;
  wire  \inst_doa_mux_b2/B0_7 ;
  wire  \inst_doa_mux_b2/B1_0 ;
  wire  \inst_doa_mux_b2/B1_1 ;
  wire  \inst_doa_mux_b2/B1_2 ;
  wire  \inst_doa_mux_b2/B1_3 ;
  wire  \inst_doa_mux_b2/B2_0 ;
  wire  \inst_doa_mux_b2/B2_1 ;
  wire \and_Naddra[15]_Naddr_o ;
  wire \and_Naddra[15]_addra_o ;
  wire \and_addra[15]_Naddra_o ;
  wire \and_addra[15]_addra[_o ;
  wire inst_doa_i0_000;
  wire inst_doa_i10_000;
  wire inst_doa_i10_001;
  wire inst_doa_i10_002;
  wire inst_doa_i11_000;
  wire inst_doa_i11_001;
  wire inst_doa_i11_002;
  wire inst_doa_i12_000;
  wire inst_doa_i12_001;
  wire inst_doa_i12_002;
  wire inst_doa_i13_000;
  wire inst_doa_i13_001;
  wire inst_doa_i14_000;
  wire inst_doa_i15_000;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i2_000;
  wire inst_doa_i2_001;
  wire inst_doa_i2_002;
  wire inst_doa_i3_000;
  wire inst_doa_i3_001;
  wire inst_doa_i3_002;
  wire inst_doa_i4_000;
  wire inst_doa_i4_001;
  wire inst_doa_i4_002;
  wire inst_doa_i5_000;
  wire inst_doa_i5_001;
  wire inst_doa_i5_002;
  wire inst_doa_i6_000;
  wire inst_doa_i6_001;
  wire inst_doa_i6_002;
  wire inst_doa_i7_000;
  wire inst_doa_i7_001;
  wire inst_doa_i7_002;
  wire inst_doa_i8_000;
  wire inst_doa_i8_001;
  wire inst_doa_i8_002;
  wire inst_doa_i9_000;
  wire inst_doa_i9_001;
  wire inst_doa_i9_002;

  assign doa[7] = doa[2];
  assign doa[6] = doa[2];
  assign doa[5] = doa[2];
  assign doa[4] = doa[2];
  assign doa[3] = doa[2];
  reg_sr_as_w1 addra_pipe_b0 (
    .clk(clka),
    .d(addra[13]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[0]));
  reg_sr_as_w1 addra_pipe_b1 (
    .clk(clka),
    .d(addra[14]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[1]));
  reg_sr_as_w1 addra_pipe_b2 (
    .clk(clka),
    .d(addra[15]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[2]));
  reg_sr_as_w1 addra_pipe_b3 (
    .clk(clka),
    .d(addra[16]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[3]));
  and \and_Naddra[15]_Naddr  (\and_Naddra[15]_Naddr_o , ~addra[15], ~addra[16]);
  and \and_Naddra[15]_addra  (\and_Naddra[15]_addra_o , ~addra[15], addra[16]);
  and \and_addra[15]_Naddra  (\and_addra[15]_Naddra_o , addra[15], ~addra[16]);
  and \and_addra[15]_addra[  (\and_addra[15]_addra[_o , addra[15], addra[16]);
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_000000_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_Naddr_o ,addra[14:13]}),
    .dia({open_n66,open_n67,open_n68,open_n69,open_n70,open_n71,open_n72,1'b0,open_n73}),
    .rsta(rsta),
    .doa({open_n88,open_n89,open_n90,open_n91,open_n92,open_n93,open_n94,open_n95,inst_doa_i0_000}));
  // address_offset=8192;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h3FFFFFFFF8000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h00007FFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000003FFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000FFFFFFFFFFFFF00000001FFFFFFFFFFFFE00),
    .INIT_18(256'hFFFFFFF800000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h00000000000000000000000000000000003FFFFFFFFFE0000000000000000FFF),
    .INIT_1A(256'h00000001FFFFFFFFC00000000000000000000000000000000000000000000000),
    .INIT_1B(256'h000000000000000000000000000000000000000007FFFFFFFF00000000000000),
    .INIT_1C(256'h000000000000000001FFFFFFFE00000000000000000000000000000000000000),
    .INIT_1D(256'h000000000000000000000000000000000000000000000000FFFFFFFF00000000),
    .INIT_1E(256'h0000000000000000000000000003FFFFFFE00000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000FFFFFFF80),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_008192_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_Naddr_o ,addra[14:13]}),
    .dia({open_n124,open_n125,open_n126,open_n127,open_n128,open_n129,open_n130,1'b0,open_n131}),
    .rsta(rsta),
    .doa({open_n146,open_n147,open_n148,open_n149,open_n150,open_n151,open_n152,open_n153,inst_doa_i1_000}));
  // address_offset=8192;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h00000000000000000000000000000000000000000FFFFFFFE000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFF000),
    .INIT_1A(256'hFFFFFFFE00000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h00000000000000000000000000000000000000000000000000FFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000),
    .INIT_1D(256'h00000000000000000000000000000000000000000000000000000000FFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000),
    .INIT_1F(256'h000000000000000000000000000000000000000000000000000000000000007F),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_008192_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_Naddr_o ,addra[14:13]}),
    .dia({open_n182,open_n183,open_n184,open_n185,open_n186,open_n187,open_n188,1'b0,open_n189}),
    .rsta(rsta),
    .doa({open_n204,open_n205,open_n206,open_n207,open_n208,open_n209,open_n210,open_n211,inst_doa_i1_001}));
  // address_offset=8192;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_008192_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_Naddr_o ,addra[14:13]}),
    .dia({open_n240,open_n241,open_n242,open_n243,open_n244,open_n245,open_n246,1'b0,open_n247}),
    .rsta(rsta),
    .doa({open_n262,open_n263,open_n264,open_n265,open_n266,open_n267,open_n268,open_n269,inst_doa_i1_002}));
  // address_offset=16384;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFC000000000000000000000000000000007FFFFFE00000000000000000000),
    .INIT_01(256'h00000000000000000000000000000000000000000000000000000000000000FF),
    .INIT_02(256'h00000FFFFFF000000000000000000000000000000000001FFFFFE00000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h000000000000FFFFFE00000000000000000000000000000000000000FFFFFE00),
    .INIT_05(256'h07FFFFE000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000FFFFFC000000000000000000000000000000000000000),
    .INIT_07(256'h00000000007FFFFC000000000000000000000000000000000000000000000000),
    .INIT_08(256'h000000000000000000000000007FFFFC00000000000000000000000000000000),
    .INIT_09(256'h00000000000000000007FFFF8000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000003FFFFC0000000000000000000000000),
    .INIT_0B(256'h00000000000000000000000000007FFFF8000000000000000000000000000000),
    .INIT_0C(256'h00000000000000000000000000000000000000003FFFFC000000000000000000),
    .INIT_0D(256'h00000000000000000000000000000000000007FFFF0000000000000000000000),
    .INIT_0E(256'h000000000000000000000000000000000000000000000001FFFFC00000000000),
    .INIT_0F(256'h00000000000000000000000000000000000000000000007FFFE0000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000FFFFC0000),
    .INIT_11(256'hFFE0000000000000000000000000000000000000000000000000000FFFF80000),
    .INIT_12(256'hFFFF00000000000000000000000000000000000000000000000000000000003F),
    .INIT_13(256'h000001FFFF000000000000000000000000000000000000000000000000000001),
    .INIT_14(256'h000000001FFFE000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000FFFF00000000000000000000000000000000000000000000000),
    .INIT_16(256'h000000000000000003FFF8000000000000000000000000000000000000000000),
    .INIT_17(256'h000000000000000000003FFF8000000000000000000000000000000000000000),
    .INIT_18(256'h000000000000000000000000007FFF0000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000001FFFC00000000000000000000000000000000),
    .INIT_1A(256'h00000000000000000000000000000000001FFFC0000000000000000000000000),
    .INIT_1B(256'h000000000000000000000000000000000007FFF0000000000000000000000000),
    .INIT_1C(256'h00000000000000000000000000000000000000000003FFF00000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000001FFF800000000000000000),
    .INIT_1E(256'h00000000000000000000000000000000000000000000000000007FFE00000000),
    .INIT_1F(256'h80000000000000000000000000000000000000000000000000FFFC0000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_016384_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_Naddr_o ,addra[14:13]}),
    .dia({open_n298,open_n299,open_n300,open_n301,open_n302,open_n303,open_n304,1'b0,open_n305}),
    .rsta(rsta),
    .doa({open_n320,open_n321,open_n322,open_n323,open_n324,open_n325,open_n326,open_n327,inst_doa_i2_000}));
  // address_offset=16384;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000),
    .INIT_05(256'hF800000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFF800000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h00000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000),
    .INIT_0A(256'h000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000),
    .INIT_0E(256'h00000000000000000000000000000000000000000000000000003FFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000),
    .INIT_10(256'h000000000000000000000000000000000000000000000000000000000003FFFF),
    .INIT_11(256'h001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE),
    .INIT_14(256'hFFFFFFFFE0000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h00000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000),
    .INIT_19(256'h00000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000),
    .INIT_1B(256'h000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000),
    .INIT_1D(256'h00000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000),
    .INIT_1F(256'h000000000000000000000000000000000000000000000000000003FFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_016384_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_Naddr_o ,addra[14:13]}),
    .dia({open_n356,open_n357,open_n358,open_n359,open_n360,open_n361,open_n362,1'b0,open_n363}),
    .rsta(rsta),
    .doa({open_n378,open_n379,open_n380,open_n381,open_n382,open_n383,open_n384,open_n385,inst_doa_i2_001}));
  // address_offset=16384;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_016384_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_Naddr_o ,addra[14:13]}),
    .dia({open_n414,open_n415,open_n416,open_n417,open_n418,open_n419,open_n420,1'b0,open_n421}),
    .rsta(rsta),
    .doa({open_n436,open_n437,open_n438,open_n439,open_n440,open_n441,open_n442,open_n443,inst_doa_i2_002}));
  // address_offset=24576;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000001FFF),
    .INIT_01(256'h000003FFE0000000000000000000000000000000000000000000000003FFF000),
    .INIT_02(256'h0FFF800000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h00000000000000FFF80000000000000000000000000000000000000000000000),
    .INIT_04(256'h000000003FFE0000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h000000007C0000000000003FFE00000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000FFF800000000006000000000000000000000000000000000),
    .INIT_07(256'h00000000000000003FE0000000000007FF800000000000000000000000000000),
    .INIT_08(256'h000000000000000000000003FFC00000000007E0000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000FFC000000000001FFE000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000FFF0000000000FFC00000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000007FF8000000000007FF8000000000000),
    .INIT_0C(256'h000000000000000000000000000000000000003FFC0000000007FF8000000000),
    .INIT_0D(256'h000000000000000000000000000000000000000003FFF000000000001FFC0000),
    .INIT_0E(256'h07FF0000000000000000000000000000000000000000007FF0000000003FFF00),
    .INIT_0F(256'h00FFFE00000000000000000000000000000000000000000001FFFE0000000000),
    .INIT_10(256'h0000000001FFC00000000000000000000000000000000000000001FFC0000000),
    .INIT_11(256'h0000000007FFFC00000000000000000000000000000000000000000000FFFFC0),
    .INIT_12(256'h003FFFF000000000007FF00000000000000000000000000000000000000007FF),
    .INIT_13(256'h00001FFC000000001FFFFC000000000000000000000000000000000000000000),
    .INIT_14(256'h00000000001FFFFC00000000003FF80000000000000000000000000000000000),
    .INIT_15(256'h0000000000003FF800000000FFFFF80000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000001FFFFF80000000000FFE00000000000000000000000000),
    .INIT_17(256'h00000000000000000000FFE000000003FFFFF000000000000000000000000000),
    .INIT_18(256'h000000000000000000000000000FFFFFC00000000003FF000000000000000000),
    .INIT_19(256'h0000000000000000000000000001FF800000000FFFFFE0000000000000000000),
    .INIT_1A(256'h000000000000000000000000000000000007FFFFF00000000000FFC000000000),
    .INIT_1B(256'h000000000000000000000000000000000007FE000000003FFFFFE00000000000),
    .INIT_1C(256'h00000000000000000000000000000000000000000003FFFFFC00000000007FE0),
    .INIT_1D(256'h00001FF800000000000000000000000000000000000FFC00000000FFFFFFC000),
    .INIT_1E(256'hFFFFC00000000000000000000000000000000000000000000003FFFFFF000000),
    .INIT_1F(256'hFFC0000000000FFC00000000000000000000000000000000003FF000000003FF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_024576_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_Naddr_o ,addra[14:13]}),
    .dia({open_n472,open_n473,open_n474,open_n475,open_n476,open_n477,open_n478,1'b0,open_n479}),
    .rsta(rsta),
    .doa({open_n494,open_n495,open_n496,open_n497,open_n498,open_n499,open_n500,open_n501,inst_doa_i3_000}));
  // address_offset=24576;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000),
    .INIT_01(256'hFFFFFC0000000000000000000000000000000000000000000000000000000FFF),
    .INIT_02(256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000),
    .INIT_04(256'h000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFF83FFFFFFFFFFFFC00000000000000000000000000000000000000000),
    .INIT_06(256'h00000000000000000007FFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFC01FFFFFFFFFFFF800000000000000000000000000000000),
    .INIT_08(256'h000000000000000000000000003FFFFFFFFFF81FFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFF003FFFFFFFFFFFE000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000FFFFFFFFFF003FFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8007FFFFFFFFFFF8000000000000000),
    .INIT_0C(256'h000000000000000000000000000000000000000003FFFFFFFFF8007FFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFFFFFFFE0000000),
    .INIT_0E(256'hF800000000000000000000000000000000000000000000000FFFFFFFFFC000FF),
    .INIT_0F(256'hFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFE00000000000000000000000000000000000000000000003FFFFFFF),
    .INIT_11(256'hFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00003F),
    .INIT_12(256'hFFC0000FFFFFFFFFFF8000000000000000000000000000000000000000000000),
    .INIT_13(256'h00000003FFFFFFFFE00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFE00003FFFFFFFFFFC0000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000007FFFFFFFF000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFE000007FFFFFFFFFF00000000000000000000000000000),
    .INIT_17(256'h00000000000000000000001FFFFFFFFC00000FFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF000003FFFFFFFFFFC00000000000000000000),
    .INIT_19(256'h0000000000000000000000000000007FFFFFFFF000001FFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000FFFFFFFFFFF000000000000),
    .INIT_1B(256'h00000000000000000000000000000000000001FFFFFFFFC000001FFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000003FFFFFFFFFF8000),
    .INIT_1D(256'hFFFFE00000000000000000000000000000000000000003FFFFFFFF0000003FFF),
    .INIT_1E(256'h00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000FFFFFF),
    .INIT_1F(256'h003FFFFFFFFFF0000000000000000000000000000000000000000FFFFFFFFC00),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_024576_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_Naddr_o ,addra[14:13]}),
    .dia({open_n530,open_n531,open_n532,open_n533,open_n534,open_n535,open_n536,1'b0,open_n537}),
    .rsta(rsta),
    .doa({open_n552,open_n553,open_n554,open_n555,open_n556,open_n557,open_n558,open_n559,inst_doa_i3_001}));
  // address_offset=24576;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_024576_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_Naddr_o ,addra[14:13]}),
    .dia({open_n588,open_n589,open_n590,open_n591,open_n592,open_n593,open_n594,1'b0,open_n595}),
    .rsta(rsta),
    .doa({open_n610,open_n611,open_n612,open_n613,open_n614,open_n615,open_n616,open_n617,inst_doa_i3_002}));
  // address_offset=32768;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000FFFFFFFC00000000000000000000000000000000000000000000003FFFF),
    .INIT_01(256'h0001FFFFFFE00000000003FF00000000000000000000000000000000007FE000),
    .INIT_02(256'h01FF800000003FFFFFFF80000000000000000000000000000000000000000000),
    .INIT_03(256'h000000000001FFFFFFF80000000001FF80000000000000000000000000000000),
    .INIT_04(256'h0000000003FF000000007FFFFFFF800000000000000000008000000000000000),
    .INIT_05(256'h00000000000000000001FFFFFFFC00000000007FC00000000000000000000000),
    .INIT_06(256'h000000000000000007FC00000001FFFFFFFF8000000000000000000080000000),
    .INIT_07(256'hC000000200000000000000000001FFFFFFFF00000000003FE000000000000000),
    .INIT_08(256'h0000000000000000000000000FF800000007FFFFFFFF00000000000000000000),
    .INIT_09(256'h00000000C000000700000000000000000001FFFFFFFF80000000000FF8000000),
    .INIT_0A(256'hFC0000000000000000000000000000003FE00000000FFFFFFFFF000000000000),
    .INIT_0B(256'h0000000000000001C000000700000000000000000001FFFFFFFFE00000000007),
    .INIT_0C(256'h00000003FE0000000000000000000000000000007FC00000003FFFFFFFFF0000),
    .INIT_0D(256'hFFFF00000000000000000001E000000F00000000000000000001FFFFFFFFF000),
    .INIT_0E(256'hFFFFFC0000000001FF000000000000000000000000000000FF800000007FFFFF),
    .INIT_0F(256'h00FFFFFFFFFF00000000000000000001E000000F00000000000000000003FFFF),
    .INIT_10(256'h0003FFFFFFFFFE00000000007F800000000000000000000000000001FF000000),
    .INIT_11(256'hFC00000003FFFFFFFFFF00000000000000000001F000000F0000000000000000),
    .INIT_12(256'h000000000003FFFFFFFFFF80000000003FC00000000000000000000000000003),
    .INIT_13(256'h00000007F800000007FFFFFFFFFF80000000000000000001F000001F00000000),
    .INIT_14(256'h00000000000000000003FFFFFFFFFFC0000000001FE000000000000000000000),
    .INIT_15(256'h000000000000000FF00000001FFFFFFFFFFF80000000000000000001F000001F),
    .INIT_16(256'hF800003F80000000000000000007FFFFFFFFFFE0000000000FF0000000000000),
    .INIT_17(256'h00000000000000000000001FE00000003FFFFFFFFFFF80000000000000000001),
    .INIT_18(256'h00000003F800003F80000000000000000007FFFFFFFFFFF80000000007F80000),
    .INIT_19(256'h03FC000000000000000000000000003FC00000007FFFFFFFFFFFC00000000000),
    .INIT_1A(256'h0000000000000003FC00003F80000000000000000007FFFFFFFFFFFC00000000),
    .INIT_1B(256'h0000000001FE000000000000000000000000007F80000000FFFFFFFFFFFFC000),
    .INIT_1C(256'hFFFFC0000000000000000003FC00007F8000000000000000000FFFFFFFFFFFFE),
    .INIT_1D(256'hFFFFFFFF0000000000FF00000000000000000000000000FF00000001FFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFE0000000000000000003FC00007F8000000000000000000FFFFF),
    .INIT_1F(256'h001FFFFFFFFFFFFF80000000007F80000000000000000000000001FE00000007),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_032768_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_Naddra_o ,addra[14:13]}),
    .dia({open_n646,open_n647,open_n648,open_n649,open_n650,open_n651,open_n652,1'b0,open_n653}),
    .rsta(rsta),
    .doa({open_n668,open_n669,open_n670,open_n671,open_n672,open_n673,open_n674,open_n675,inst_doa_i4_000}));
  // address_offset=32768;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFF00000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000),
    .INIT_01(256'hFFFE0000001FFFFFFFFFFC000000000000000000000000000000000000001FFF),
    .INIT_02(256'h00007FFFFFFFC00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFE00000007FFFFFFFFFE0000000000000000000000000000000000),
    .INIT_04(256'h000000000000FFFFFFFF800000007FFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFE00000003FFFFFFFFFF80000000000000000000000000),
    .INIT_06(256'h00000000000000000003FFFFFFFE000000007FFFFFFFFFFFFFFFFFFF7FFFFFFF),
    .INIT_07(256'h3FFFFFFDFFFFFFFFFFFFFFFFFFFE00000000FFFFFFFFFFC00000000000000000),
    .INIT_08(256'h0000000000000000000000000007FFFFFFF800000000FFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFF3FFFFFF8FFFFFFFFFFFFFFFFFFFE000000007FFFFFFFFFF000000000),
    .INIT_0A(256'h00000000000000000000000000000000001FFFFFFFF000000000FFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFE3FFFFFF8FFFFFFFFFFFFFFFFFFFE000000001FFFFFFFFFF8),
    .INIT_0C(256'hFFFFFFFC00000000000000000000000000000000003FFFFFFFC000000000FFFF),
    .INIT_0D(256'h0000FFFFFFFFFFFFFFFFFFFE1FFFFFF0FFFFFFFFFFFFFFFFFFFE000000000FFF),
    .INIT_0E(256'h000003FFFFFFFFFE00000000000000000000000000000000007FFFFFFF800000),
    .INIT_0F(256'hFF0000000000FFFFFFFFFFFFFFFFFFFE1FFFFFF0FFFFFFFFFFFFFFFFFFFC0000),
    .INIT_10(256'hFFFC0000000001FFFFFFFFFF8000000000000000000000000000000000FFFFFF),
    .INIT_11(256'h03FFFFFFFC0000000000FFFFFFFFFFFFFFFFFFFE0FFFFFF0FFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFC00000000007FFFFFFFFFC0000000000000000000000000000000),
    .INIT_13(256'h0000000007FFFFFFF800000000007FFFFFFFFFFFFFFFFFFE0FFFFFE0FFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFC00000000003FFFFFFFFFE00000000000000000000000),
    .INIT_15(256'h00000000000000000FFFFFFFE000000000007FFFFFFFFFFFFFFFFFFE0FFFFFE0),
    .INIT_16(256'h07FFFFC07FFFFFFFFFFFFFFFFFF800000000001FFFFFFFFFF000000000000000),
    .INIT_17(256'h0000000000000000000000001FFFFFFFC000000000007FFFFFFFFFFFFFFFFFFE),
    .INIT_18(256'hFFFFFFFC07FFFFC07FFFFFFFFFFFFFFFFFF8000000000007FFFFFFFFF8000000),
    .INIT_19(256'hFC0000000000000000000000000000003FFFFFFF8000000000003FFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFC03FFFFC07FFFFFFFFFFFFFFFFFF8000000000003FFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFE0000000000000000000000000000007FFFFFFF0000000000003FFF),
    .INIT_1C(256'h00003FFFFFFFFFFFFFFFFFFC03FFFF807FFFFFFFFFFFFFFFFFF0000000000001),
    .INIT_1D(256'h00000000FFFFFFFFFF000000000000000000000000000000FFFFFFFE00000000),
    .INIT_1E(256'h0000000000001FFFFFFFFFFFFFFFFFFC03FFFF807FFFFFFFFFFFFFFFFFF00000),
    .INIT_1F(256'hFFE00000000000007FFFFFFFFF800000000000000000000000000001FFFFFFF8),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_032768_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_Naddra_o ,addra[14:13]}),
    .dia({open_n704,open_n705,open_n706,open_n707,open_n708,open_n709,open_n710,1'b0,open_n711}),
    .rsta(rsta),
    .doa({open_n726,open_n727,open_n728,open_n729,open_n730,open_n731,open_n732,open_n733,inst_doa_i4_001}));
  // address_offset=32768;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_032768_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_Naddra_o ,addra[14:13]}),
    .dia({open_n762,open_n763,open_n764,open_n765,open_n766,open_n767,open_n768,1'b0,open_n769}),
    .rsta(rsta),
    .doa({open_n784,open_n785,open_n786,open_n787,open_n788,open_n789,open_n790,open_n791,inst_doa_i4_002}));
  // address_offset=40960;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000FFFFFFFFFFFFFE0000000000000000003FE0000FF8000000000000000),
    .INIT_01(256'h00000000001FFFFFFFFFFFFFE0000000003F80000000000000000000000003FC),
    .INIT_02(256'h000003F80000001FFFFFFFFFFFFFF0000000000000000003FE0000FF80000000),
    .INIT_03(256'h8000000000000000003FFFFFFFFFFFFFF0000000001FC0000000000000000000),
    .INIT_04(256'h00000000000007F00000003FFFFFFFFFFFFFF8000000000000000003FE0000FF),
    .INIT_05(256'hFF0001FF8000000000000000007FFFFFFFFFFFFFF8000000000FE00000000000),
    .INIT_06(256'h000000000000000000000FE00000007FFFFFFFFFFFFFF8000000000000000007),
    .INIT_07(256'h00000007FF0001FF8000000000000000007FFFFFFFFFFFFFFC0000000007F000),
    .INIT_08(256'h0007F000000000000000000000001FC0000000FFFFFFFFFFFFFFFC0000000000),
    .INIT_09(256'h0000000000000007FF8001FFC00000000000000000FFFFFFFFFFFFFFFE000000),
    .INIT_0A(256'hFF0000000003F800000000000000000000001FC0000001FFFFFFFFFFFFFFFF00),
    .INIT_0B(256'hFFFFFF000000000000000007FF8003FFC00000000000000001FFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFF8000000001FC00000000000000000000003F80000003FFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFF800000000000000007FFFFFFFFC00000000000000003FFFFFF),
    .INIT_0E(256'h07FFFFFFFFFFFFFFFFC000000000FC00000000000000000000007F00000007FF),
    .INIT_0F(256'h00000FFFFFFFFFFFFFFFFFC00000000000000007FFFFFFFFC000000000000000),
    .INIT_10(256'h000000000FFFFFFFFFFFFFFFFFE000000000FE00000000000000000000007E00),
    .INIT_11(256'h0000FE0000001FFFFFFFFFFFFFFFFFF00000000000000007FFFFFFFFC0000000),
    .INIT_12(256'hE0000000000000001FFFFFFFFFFFFFFFFFF0000000007F000000000000000000),
    .INIT_13(256'h000000000001FC0000003FFFFFFFFFFFFFFFFFF8000000000000000FFFFFFFFF),
    .INIT_14(256'hFFFFFFFFE0000000000000007FFFFFFFFFFFFFFFFFF8000000003F0000000000),
    .INIT_15(256'h00000000000000000001F80000007FFFFFFFFFFFFFFFFFFE000000000000000F),
    .INIT_16(256'h0000000FFFFFFFFFE000000000000000FFFFFFFFFFFFFFFFFFFC000000003F80),
    .INIT_17(256'h00001F8000000000000000000003F8000000FFFFFFFFFFFFFFFFFFFF00000000),
    .INIT_18(256'hC00000000000000FFFFFFFFFE000000000000003FFFFFFFFFFFFFFFFFFFE0000),
    .INIT_19(256'hFFFF000000000FC000000000000000000003F0000001FFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFF00000000000000FFFFFFFFFE00000000000000FFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFF000000000FC000000000000000000007E0000003FFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFC0000000000001FFFFFFFFFF00000000000001FFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFF8000000007E000000000000000000007E0000003FFFF),
    .INIT_1E(256'h0007FFFFFFFFFFFFFFFFFFFFFF0000000000001FFFFFFFFFF00000000000007F),
    .INIT_1F(256'h000003FFFFFFFFFFFFFFFFFFFFFFC000000007E00000000000000000000FC000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_040960_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_Naddra_o ,addra[14:13]}),
    .dia({open_n820,open_n821,open_n822,open_n823,open_n824,open_n825,open_n826,1'b0,open_n827}),
    .rsta(rsta),
    .doa({open_n842,open_n843,open_n844,open_n845,open_n846,open_n847,open_n848,open_n849,inst_doa_i5_000}));
  // address_offset=40960;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFF00000000000001FFFFFFFFFFFFFFFFFFC01FFFF007FFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFE00000000000001FFFFFFFFFC00000000000000000000000000003),
    .INIT_02(256'h00000007FFFFFFE00000000000000FFFFFFFFFFFFFFFFFFC01FFFF007FFFFFFF),
    .INIT_03(256'h7FFFFFFFFFFFFFFFFFC00000000000000FFFFFFFFFE000000000000000000000),
    .INIT_04(256'h000000000000000FFFFFFFC000000000000007FFFFFFFFFFFFFFFFFC01FFFF00),
    .INIT_05(256'h00FFFE007FFFFFFFFFFFFFFFFF8000000000000007FFFFFFFFF0000000000000),
    .INIT_06(256'h00000000000000000000001FFFFFFF8000000000000007FFFFFFFFFFFFFFFFF8),
    .INIT_07(256'hFFFFFFF800FFFE007FFFFFFFFFFFFFFFFF8000000000000003FFFFFFFFF80000),
    .INIT_08(256'hFFF8000000000000000000000000003FFFFFFF0000000000000003FFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFF8007FFE003FFFFFFFFFFFFFFFFF0000000000000001FFFFFF),
    .INIT_0A(256'h00FFFFFFFFFC000000000000000000000000003FFFFFFE0000000000000000FF),
    .INIT_0B(256'h000000FFFFFFFFFFFFFFFFF8007FFC003FFFFFFFFFFFFFFFFE00000000000000),
    .INIT_0C(256'h00000000007FFFFFFFFE000000000000000000000000007FFFFFFC0000000000),
    .INIT_0D(256'h000000000000007FFFFFFFFFFFFFFFF8000000003FFFFFFFFFFFFFFFFC000000),
    .INIT_0E(256'hF800000000000000003FFFFFFFFF00000000000000000000000000FFFFFFF800),
    .INIT_0F(256'hFFFFF000000000000000003FFFFFFFFFFFFFFFF8000000003FFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFF000000000000000001FFFFFFFFF00000000000000000000000001FF),
    .INIT_11(256'h000001FFFFFFE000000000000000000FFFFFFFFFFFFFFFF8000000003FFFFFFF),
    .INIT_12(256'h1FFFFFFFFFFFFFFFE000000000000000000FFFFFFFFF80000000000000000000),
    .INIT_13(256'h00000000000003FFFFFFC0000000000000000007FFFFFFFFFFFFFFF000000000),
    .INIT_14(256'h000000001FFFFFFFFFFFFFFF80000000000000000007FFFFFFFFC00000000000),
    .INIT_15(256'h0000000000000000000007FFFFFF80000000000000000001FFFFFFFFFFFFFFF0),
    .INIT_16(256'hFFFFFFF0000000001FFFFFFFFFFFFFFF00000000000000000003FFFFFFFFC000),
    .INIT_17(256'hFFFFE0000000000000000000000007FFFFFF00000000000000000000FFFFFFFF),
    .INIT_18(256'h3FFFFFFFFFFFFFF0000000001FFFFFFFFFFFFFFC00000000000000000001FFFF),
    .INIT_19(256'h0000FFFFFFFFF000000000000000000000000FFFFFFE00000000000000000000),
    .INIT_1A(256'h000000000FFFFFFFFFFFFFF0000000001FFFFFFFFFFFFFF00000000000000000),
    .INIT_1B(256'h000000000000FFFFFFFFF000000000000000000000001FFFFFFC000000000000),
    .INIT_1C(256'h000000000000000003FFFFFFFFFFFFE0000000000FFFFFFFFFFFFFE000000000),
    .INIT_1D(256'h000000000000000000007FFFFFFFF800000000000000000000001FFFFFFC0000),
    .INIT_1E(256'hFFF80000000000000000000000FFFFFFFFFFFFE0000000000FFFFFFFFFFFFF80),
    .INIT_1F(256'hFFFFFC00000000000000000000003FFFFFFFF800000000000000000000003FFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_040960_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_Naddra_o ,addra[14:13]}),
    .dia({open_n878,open_n879,open_n880,open_n881,open_n882,open_n883,open_n884,1'b0,open_n885}),
    .rsta(rsta),
    .doa({open_n900,open_n901,open_n902,open_n903,open_n904,open_n905,open_n906,open_n907,inst_doa_i5_001}));
  // address_offset=40960;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_040960_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_Naddra_o ,addra[14:13]}),
    .dia({open_n936,open_n937,open_n938,open_n939,open_n940,open_n941,open_n942,1'b0,open_n943}),
    .rsta(rsta),
    .doa({open_n958,open_n959,open_n960,open_n961,open_n962,open_n963,open_n964,open_n965,inst_doa_i5_002}));
  // address_offset=49152;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000FC000000FFFFFFFFFFFFFFFFFFFFFFFC000000000001FFFFFFFFFF0000000),
    .INIT_01(256'hF000000000001FFFFFFFFFFFFFFFFFFFFFFFE000000003F00000000000000000),
    .INIT_02(256'h00000000001F8000001FFFFFFFFFFFFFFFFFFFFFFFF800000000001FFFFFFFFF),
    .INIT_03(256'hFFFFFFFFF80000000000FFFFFFFFFFFFFFFFFFFFFFFFF000000003F000000000),
    .INIT_04(256'h0000000000000000001F8000003FFFFFFFFFFFFFFFFFFFFFFFFF00000000003F),
    .INIT_05(256'h0000003FFFFFFFFFF80000000007FFFFFFFFFFFFFFFFFFFFFFFFF000000001F0),
    .INIT_06(256'h000001F80000000000000000001F0000003FFFFFFFFFFFFFFFFFFFFFFFFFE000),
    .INIT_07(256'hFFFFFE000000003FFFFFFFFFF8000000007FFFFFFFFFFFFFFFFFFFFFFFFFF800),
    .INIT_08(256'hFFFFFC00000001F80000000000000000003F0000007FFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFE00000003FFFFFFFFFFC0000000FFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFE00000000F80000000000000000003F000000FFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFF8000007FFFFFFFFFFC00000FFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFE00000000FC0000000000000000003E000000FFFFFF),
    .INIT_0D(256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000FFFFFFFFFFFE00FFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000FC0000000000000000007E0000),
    .INIT_0F(256'h007E000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000007C0000000000000000),
    .INIT_11(256'h00000000007C000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000007E00000000),
    .INIT_13(256'h000000000000000000FC000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000007E),
    .INIT_15(256'h0000003E000000000000000000FC000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0),
    .INIT_17(256'hFFFFFFE00000003E000000000000000000F800000FFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFE00000003E000000000000000000F800001FFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFF00000003E000000000000000000F800001FFFFFFF),
    .INIT_1C(256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000003F000000000000000000F80000),
    .INIT_1E(256'h01F800003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000003F0000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_049152_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_Naddra_o ,addra[14:13]}),
    .dia({open_n994,open_n995,open_n996,open_n997,open_n998,open_n999,open_n1000,1'b0,open_n1001}),
    .rsta(rsta),
    .doa({open_n1016,open_n1017,open_n1018,open_n1019,open_n1020,open_n1021,open_n1022,open_n1023,inst_doa_i6_000}));
  // address_offset=49152;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00003FFFFFF000000000000000000000003FFFFFFFFFFFE0000000000FFFFFFF),
    .INIT_01(256'h0FFFFFFFFFFFE000000000000000000000001FFFFFFFFC000000000000000000),
    .INIT_02(256'h0000000000007FFFFFE0000000000000000000000007FFFFFFFFFFE000000000),
    .INIT_03(256'h0000000007FFFFFFFFFF0000000000000000000000000FFFFFFFFC0000000000),
    .INIT_04(256'h000000000000000000007FFFFFC0000000000000000000000000FFFFFFFFFFC0),
    .INIT_05(256'hFFFFFFC00000000007FFFFFFFFF80000000000000000000000000FFFFFFFFE00),
    .INIT_06(256'hFFFFFE0000000000000000000000FFFFFFC00000000000000000000000001FFF),
    .INIT_07(256'h000001FFFFFFFFC00000000007FFFFFFFF8000000000000000000000000007FF),
    .INIT_08(256'h000003FFFFFFFE0000000000000000000000FFFFFF8000000000000000000000),
    .INIT_09(256'h000000000000001FFFFFFFC00000000003FFFFFFF00000000000000000000000),
    .INIT_0A(256'h00000000000001FFFFFFFF0000000000000000000000FFFFFF00000000000000),
    .INIT_0B(256'h0000000000000000000000007FFFFF800000000003FFFFF00000000000000000),
    .INIT_0C(256'h0000000000000000000001FFFFFFFF0000000000000000000001FFFFFF000000),
    .INIT_0D(256'hFE000000000000000000000000000000001FFF000000000001FF000000000000),
    .INIT_0E(256'h000000000000000000000000000000FFFFFFFF0000000000000000000001FFFF),
    .INIT_0F(256'h0001FFFFFC000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h00000000000000000000000000000000000000FFFFFFFF800000000000000000),
    .INIT_11(256'h000000000003FFFFFC0000000000000000000000000000000000000000000000),
    .INIT_12(256'h00000000000000000000000000000000000000000000007FFFFFFF8000000000),
    .INIT_13(256'h00000000000000000003FFFFF800000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000003FFFFFFF80),
    .INIT_15(256'hFFFFFFC000000000000000000003FFFFF8000000000000000000000000000000),
    .INIT_16(256'h000000000000000000000000000000000000000000000000000000000000003F),
    .INIT_17(256'h0000001FFFFFFFC000000000000000000007FFFFF00000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h000000000000001FFFFFFFC000000000000000000007FFFFE000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h00000000000000000000000FFFFFFFC000000000000000000007FFFFE0000000),
    .INIT_1C(256'hC000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000FFFFFFFC000000000000000000007FFFF),
    .INIT_1E(256'h0007FFFFC0000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000007FFFFFFC00000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_049152_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_Naddra_o ,addra[14:13]}),
    .dia({open_n1052,open_n1053,open_n1054,open_n1055,open_n1056,open_n1057,open_n1058,1'b0,open_n1059}),
    .rsta(rsta),
    .doa({open_n1074,open_n1075,open_n1076,open_n1077,open_n1078,open_n1079,open_n1080,open_n1081,inst_doa_i6_001}));
  // address_offset=49152;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_049152_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_Naddra_o ,addra[14:13]}),
    .dia({open_n1110,open_n1111,open_n1112,open_n1113,open_n1114,open_n1115,open_n1116,1'b0,open_n1117}),
    .rsta(rsta),
    .doa({open_n1132,open_n1133,open_n1134,open_n1135,open_n1136,open_n1137,open_n1138,open_n1139,inst_doa_i6_002}));
  // address_offset=57344;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000001F800007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000001F00000000),
    .INIT_02(256'h000000000000000001F000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000001F),
    .INIT_04(256'h0000001F000000000000000001F000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC),
    .INIT_06(256'hFFFFFFFE0000001F000000000000000001F00000FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFE0000001F000000000000000001F00000FFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFE0000001F000000000000000001F00001FFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF07FFFFFFFFFFC1FFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000001F000000000000000001F00001),
    .INIT_0D(256'h01F00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0FFFFFFFFFFFE07FFFF),
    .INIT_0E(256'hFF01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000001F0000000000000000),
    .INIT_0F(256'h0000000001F00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00FFFFFFFFFF),
    .INIT_10(256'hFFEFFFFFFF007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000001F00000000),
    .INIT_11(256'h000000000000000001F00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC01FF),
    .INIT_12(256'hFFF801FFFFE7EFFFFF003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000001F),
    .INIT_13(256'h8000003F000000000000000001F00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFE001FFFFE7CFFFFF000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFF8000003F000000000000000001F80007FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFC000FFFFE7CFFFFE0007FFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFC000003E000000000000000001F80007FFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFE38FFFFE0003FFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFC000003E000000000000000000F80007FFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFE18FFFFC0001FFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000003E000000000000000000F80007),
    .INIT_1C(256'h00F80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001FFFC007FFF80000FF),
    .INIT_1D(256'hE000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000003E0000000000000000),
    .INIT_1E(256'h0000000000F8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000FFFC007FF),
    .INIT_1F(256'hFFC007FF8000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000007E00000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_057344_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_Naddra_o ,addra[14:13]}),
    .dia({open_n1168,open_n1169,open_n1170,open_n1171,open_n1172,open_n1173,open_n1174,1'b0,open_n1175}),
    .rsta(rsta),
    .doa({open_n1190,open_n1191,open_n1192,open_n1193,open_n1194,open_n1195,open_n1196,open_n1197,inst_doa_i7_000}));
  // address_offset=57344;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000000000007FFFF800000000000000000000000000000000000000000000000),
    .INIT_01(256'h000000000000000000000000000000000000000000000007FFFFFFE000000000),
    .INIT_02(256'h0000000000000000000FFFFF8000000000000000000000000000000000000000),
    .INIT_03(256'h00000000000000000000000000000000000000000000000000000003FFFFFFE0),
    .INIT_04(256'hFFFFFFE00000000000000000000FFFFF80000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000003),
    .INIT_06(256'h00000001FFFFFFE00000000000000000000FFFFF000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000001FFFFFFE00000000000000000000FFFFF0000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h000000000000000000000001FFFFFFE00000000000000000000FFFFE00000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h00000000000000000000000000000000FFFFFFE00000000000000000000FFFFE),
    .INIT_0D(256'h000FFFFE00000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000FFFFFFE00000000000000000),
    .INIT_0F(256'h00000000000FFFFC000000000000000000000000000000000000000000000000),
    .INIT_10(256'h000000000000000000000000000000000000000000000000FFFFFFE000000000),
    .INIT_11(256'h0000000000000000000FFFFC0000000000000000000000000000000000000000),
    .INIT_12(256'h000000000000000000000000000000000000000000000000000000007FFFFFE0),
    .INIT_13(256'h7FFFFFC00000000000000000000FFFFC00000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h000000007FFFFFC000000000000000000007FFF8000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h00000000000000003FFFFFC000000000000000000007FFF80000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000003FFFFFC000000000000000000007FFF800000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h000000000000000000000000000000003FFFFFC000000000000000000007FFF8),
    .INIT_1C(256'h0007FFF800000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h00000000000000000000000000000000000000001FFFFFC00000000000000000),
    .INIT_1E(256'h000000000007FFF0000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000001FFFFF8000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_057344_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_Naddra_o ,addra[14:13]}),
    .dia({open_n1226,open_n1227,open_n1228,open_n1229,open_n1230,open_n1231,open_n1232,1'b0,open_n1233}),
    .rsta(rsta),
    .doa({open_n1248,open_n1249,open_n1250,open_n1251,open_n1252,open_n1253,open_n1254,open_n1255,inst_doa_i7_001}));
  // address_offset=57344;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_057344_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_Naddra_o ,addra[14:13]}),
    .dia({open_n1284,open_n1285,open_n1286,open_n1287,open_n1288,open_n1289,open_n1290,1'b0,open_n1291}),
    .rsta(rsta),
    .doa({open_n1306,open_n1307,open_n1308,open_n1309,open_n1310,open_n1311,open_n1312,open_n1313,inst_doa_i7_002}));
  // address_offset=65536;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000000000000000000FC000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000001),
    .INIT_01(256'hF00000003FC007F80000003FFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFE000007E),
    .INIT_02(256'hE000007C000000000000000000FC000FFFFFFC0003FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFF0000000000000000000001FFFFFFFFFFFFFFFFFFFFF000000007FFF),
    .INIT_04(256'h000001FFE00000FC0000000000000000007C000FFFFC00000001FFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFE0000000000000000000000FFFFFFFFFFFFFFFFFFFC00000),
    .INIT_06(256'hFC0000000000000FF00000FC0000000000000000007E000FFE000000000007FF),
    .INIT_07(256'h0000007FFFFFFFFFFFFFFFFFE0000000000000000000000FFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFE000000000000000F00000F80000000000000000007E000FE0000000),
    .INIT_09(256'h000000000000000FFFFFFFFFFFFFFFFFC00000000000000000000007FFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFF0000000000000000000001F80000000000000000003E000F),
    .INIT_0B(256'h003F00000000000000000001FFFFFFFFFFFFFFFFC00000000000000000000007),
    .INIT_0C(256'h00000007FFFFFFFFFFFFFFFC0000000000000000000001F80000000000000000),
    .INIT_0D(256'h00000000003F000000000000000000007FFFFFFFFFFFFFFFC000000000000000),
    .INIT_0E(256'h0000000000000003FFFFFFFFFFFFFFF00000000000000000000001F000000000),
    .INIT_0F(256'h0000000000000000001F000000000000000000001FFFFFFFFFFFFFFF80000000),
    .INIT_10(256'h800000000000000000000003FFFFFFFFFFFFFFC00000000000000000000003F0),
    .INIT_11(256'h000003F00000000000000000001F8000000000000000000007FFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFF9FFF8000000000000003FFF3FFFFFFFFFFFFFF800000000000000000),
    .INIT_13(256'h00000000000007E00000000000000000001F8000000000000000000001FFFFFF),
    .INIT_14(256'h00FFFFFFFFFFFFFFFFFFF00000000000000FFFFFFFFFFFFFFFFFFF0000000000),
    .INIT_15(256'h0000000000000000000007E00000000000000000000FC0000000000000000000),
    .INIT_16(256'h00000000003FFFFFFFFFFFFFFFFFF80000000000003FFFFFFFFFFFFFFFFFFE00),
    .INIT_17(256'hFFFFF800000000000000000000000FC00000000000000000000FC00000000000),
    .INIT_18(256'h0000000000000000001FFFFFFFFFFFFFFFFFFC0000000000007FFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFF000000000000000000000000FC000000000000000000007E000),
    .INIT_1A(256'h0007E0000000000000000000000FFFFFFFFFFFFFFFFFFE0000000000007FFFFF),
    .INIT_1B(256'h00FFFFFFFFFFFFFFFFFFF000000000000000000000001F800000000000000000),
    .INIT_1C(256'h000000000003F00000000000000000000007FFFFFFFFFFFFFFFFFE0000000000),
    .INIT_1D(256'hE0000007F0FFFFFFFFFFFFFFFFFFE000000000000000000000003F8000000000),
    .INIT_1E(256'h00000000000000000003F80000000000000000000003FFFFFFFFFFFFFFFFFE1F),
    .INIT_1F(256'hFFFFFE7FF800003FFCFFFFFFFFFFFFFFFFFFC000000000000000000000003F00),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_065536_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_addra_o ,addra[14:13]}),
    .dia({open_n1342,open_n1343,open_n1344,open_n1345,open_n1346,open_n1347,open_n1348,1'b0,open_n1349}),
    .rsta(rsta),
    .doa({open_n1364,open_n1365,open_n1366,open_n1367,open_n1368,open_n1369,open_n1370,open_n1371,inst_doa_i8_000}));
  // address_offset=65536;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000003FFF00000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000001FFFF0000001FFFFF80),
    .INIT_02(256'h1FFFFF8000000000000000000003FFF0000003FFFC0000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000FFFFFFFF8000),
    .INIT_04(256'hFFFFFE001FFFFF0000000000000000000003FFF00003FFFFFFFE000000000000),
    .INIT_05(256'h00000000000000000000000000000000000000000000000000000000003FFFFF),
    .INIT_06(256'h03FFFFFFFFFFFFF00FFFFF0000000000000000000001FFF001FFFFFFFFFFF800),
    .INIT_07(256'hFFFFFF8000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h000000001FFFFFFFFFFFFFFF0FFFFF0000000000000000000001FFF01FFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFE0000000000000000000001FFF0),
    .INIT_0B(256'h0000FFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000),
    .INIT_0C(256'h000000000000000000000003FFFFFFFFFFFFFFFFFFFFFE000000000000000000),
    .INIT_0D(256'h000000000000FFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFE0000000000),
    .INIT_0F(256'h00000000000000000000FFFFFFFFFFFFFFFFFFFFE00000000000000000000000),
    .INIT_10(256'h000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFC00),
    .INIT_11(256'hFFFFFC00000000000000000000007FFFFFFFFFFFFFFFFFFFF800000000000000),
    .INIT_12(256'h00000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFF800000000000000000000007FFFFFFFFFFFFFFFFFFFFE000000),
    .INIT_14(256'hFF0000000000000000000000000000000000000000000000000000FFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFF800000000000000000000003FFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFC000000000000000000000000000000000000000000000000001FF),
    .INIT_17(256'h000007FFFFFFFFFFFFFFFFFFFFFFF000000000000000000000003FFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000001FFF),
    .INIT_1A(256'h00001FFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000),
    .INIT_1B(256'h000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000),
    .INIT_1C(256'h0000000000000FFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000),
    .INIT_1D(256'h00000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFC00000000000),
    .INIT_1E(256'h0000000000000000000007FFFFFFFFFFFFFFFFFFFFFC00000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFC000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_065536_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_addra_o ,addra[14:13]}),
    .dia({open_n1400,open_n1401,open_n1402,open_n1403,open_n1404,open_n1405,open_n1406,1'b0,open_n1407}),
    .rsta(rsta),
    .doa({open_n1422,open_n1423,open_n1424,open_n1425,open_n1426,open_n1427,open_n1428,open_n1429,inst_doa_i8_001}));
  // address_offset=65536;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_065536_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_addra_o ,addra[14:13]}),
    .dia({open_n1458,open_n1459,open_n1460,open_n1461,open_n1462,open_n1463,open_n1464,1'b0,open_n1465}),
    .rsta(rsta),
    .doa({open_n1480,open_n1481,open_n1482,open_n1483,open_n1484,open_n1485,open_n1486,open_n1487,inst_doa_i8_002}));
  // address_offset=73728;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00007F0000000000000000000001F80000000000000000000001FFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFF80000000000000000000),
    .INIT_02(256'h000000000000FE0000000000000000000001FC0000000000000000000001FFFF),
    .INIT_03(256'h0000FFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFF800000000000),
    .INIT_04(256'h00000000000000000000FC0000000000000000000000FE000000000000000000),
    .INIT_05(256'h000000000000FFFFFFFFFFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFF0000),
    .INIT_06(256'hFFFF000000000000000000000001FC00000000000000000000007E0000000000),
    .INIT_07(256'h000000000000000000007FFFFFFFFFFFFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFE000000000000000000000003F800000000000000000000007F00),
    .INIT_09(256'h00003F80000000000000000000007FFFFFFFFFFFFFFFFFFFFFF01FFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFE000000000000000000000007F0000000000000000000),
    .INIT_0B(256'h0000000000001FC0000000000000000000007FFFFFFFFFFFFFFFFFFFFFF01FFF),
    .INIT_0C(256'hFFF83FFFFFFFFFFFFFFFFFFFFFFE000000000000000000000007F00000000000),
    .INIT_0D(256'h000000000000000000001FC0000000000000000000007FFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000FE000),
    .INIT_0F(256'h001FC000000000000000000000000FE0000000000000000000007FFFFFFFFFFF),
    .INIT_10(256'hFC0001FFFFFFFFFFFFFE7FFFFFFFFFFFFF8000FFFFFC00000000000000000000),
    .INIT_11(256'h00000000003F80000000000000000000000007F0000000000000000000003FFF),
    .INIT_12(256'h00003FFFC000000FFFFFFFFFFFFEFFFFFFFFFFFFF0000007FFFC000000000000),
    .INIT_13(256'h0000000000000000007F80000000000000000000000003F80000000000000000),
    .INIT_14(256'h0000000000003FFE00000001FFFFFFFFFFFFFFFFFFFFFFFF80000000FFFC0000),
    .INIT_15(256'h3FFC0000000000000000000000FF00000000000000000000000003FC00000000),
    .INIT_16(256'h000000000000000000003FF0000000003FFFFFFFFFFFFFFFFFFFFFFC00000000),
    .INIT_17(256'h0000000007FC0000000000000000000001FE00000000000000000000000001FE),
    .INIT_18(256'h000000FF000000000000000000007FC0000000000FFFFFFFFFFFFFFFFFFFFFE0),
    .INIT_19(256'hFFFFFF800000000003FC0000000000000000000003FC00000000000000000000),
    .INIT_1A(256'h000000000000007F800000000000000000007F000000000003FFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFE000000000000FC0000000000000000000007F8000000000000),
    .INIT_1C(256'h00000000000000000000003FC00000000000000000007C0000000000007FFFFF),
    .INIT_1D(256'h003FFFFFFFFFFFFFFFFFF80000000000007C000000000000000000000FF00000),
    .INIT_1E(256'h1FE0000000000000000000000000001FE0000000000000000000780000000000),
    .INIT_1F(256'h00000000000FFFFFFFFFFFFFFFFFE00000000000001800000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_073728_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_addra_o ,addra[14:13]}),
    .dia({open_n1516,open_n1517,open_n1518,open_n1519,open_n1520,open_n1521,open_n1522,1'b0,open_n1523}),
    .rsta(rsta),
    .doa({open_n1538,open_n1539,open_n1540,open_n1541,open_n1542,open_n1543,open_n1544,open_n1545,inst_doa_i9_000}));
  // address_offset=73728;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFF80000000000000000000000007FFFFFFFFFFFFFFFFFFFFFE000000000000),
    .INIT_01(256'h000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFF00000000000000000000000003FFFFFFFFFFFFFFFFFFFFFE0000),
    .INIT_03(256'hFFFF0000000000000000000000000000000000000000000000007FFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFF00000000000000000000000001FFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFF000000000000000000000000000000000000000000000000FFFF),
    .INIT_06(256'h0000FFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000001FFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000),
    .INIT_08(256'h000000000001FFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000FF),
    .INIT_09(256'h0000007FFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000),
    .INIT_0A(256'h00000000000000000001FFFFFFFFFFFFFFFFFFFFFFF800000000000000000000),
    .INIT_0B(256'h000000000000003FFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF8000000000000),
    .INIT_0D(256'h00000000000000000000003FFFFFFFFFFFFFFFFFFFFF80000000000000000000),
    .INIT_0E(256'h000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF00000),
    .INIT_0F(256'hFFE0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFF800000000000),
    .INIT_10(256'h03FFFE00000000000000000000000000007FFF000003FFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFC0000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFC000),
    .INIT_12(256'hFFFFC0003FFFFFF00000000000000000000000000FFFFFF80003FFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFF800000000000000000000000000007FFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFC001FFFFFFFE0000000000000000000000007FFFFFFF0003FFFF),
    .INIT_15(256'hC003FFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000003FFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFC00FFFFFFFFFC00000000000000000000003FFFFFFFF),
    .INIT_17(256'hFFFFFFFFF803FFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000001),
    .INIT_18(256'h00000000FFFFFFFFFFFFFFFFFFFF803FFFFFFFFFF0000000000000000000001F),
    .INIT_19(256'h0000007FFFFFFFFFFC03FFFFFFFFFFFFFFFFFFFFFC0000000000000000000000),
    .INIT_1A(256'h00000000000000007FFFFFFFFFFFFFFFFFFF80FFFFFFFFFFFC00000000000000),
    .INIT_1B(256'h00000000000001FFFFFFFFFFFF03FFFFFFFFFFFFFFFFFFFFF800000000000000),
    .INIT_1C(256'h0000000000000000000000003FFFFFFFFFFFFFFFFFFF83FFFFFFFFFFFF800000),
    .INIT_1D(256'hFFC0000000000000000007FFFFFFFFFFFF83FFFFFFFFFFFFFFFFFFFFF0000000),
    .INIT_1E(256'hE00000000000000000000000000000001FFFFFFFFFFFFFFFFFFF87FFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFF000000000000000001FFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_073728_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_addra_o ,addra[14:13]}),
    .dia({open_n1574,open_n1575,open_n1576,open_n1577,open_n1578,open_n1579,open_n1580,1'b0,open_n1581}),
    .rsta(rsta),
    .doa({open_n1596,open_n1597,open_n1598,open_n1599,open_n1600,open_n1601,open_n1602,open_n1603,inst_doa_i9_001}));
  // address_offset=73728;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_073728_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_addra_o ,addra[14:13]}),
    .dia({open_n1632,open_n1633,open_n1634,open_n1635,open_n1636,open_n1637,open_n1638,1'b0,open_n1639}),
    .rsta(rsta),
    .doa({open_n1654,open_n1655,open_n1656,open_n1657,open_n1658,open_n1659,open_n1660,open_n1661,inst_doa_i9_002}));
  // address_offset=81920;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000000003FC0000000000000000000000000000FF00000000000000000007000),
    .INIT_01(256'h00004000000000000003FFFFFFFFFFFFFFFFC000000000000000000000000000),
    .INIT_02(256'h00000000000000007F800000000000000000000000000007F800000000000000),
    .INIT_03(256'h0000000000000000000000000001FFFFFFFFFFFFFFFF00000000000000000000),
    .INIT_04(256'h000000000000000000000001FF000000000000000000000000000003FC000000),
    .INIT_05(256'hFF00000000000000000000000000000000007FFFFFFFFFFFFFFC000000000000),
    .INIT_06(256'h00000000000000000000000000000003FE000000000000000000000000000001),
    .INIT_07(256'h00000000FF80000000000000000000000000000000003FFFFFFFFFFFFFF80000),
    .INIT_08(256'hFFE0000000000000000000000000000000000007FC0000000000000000000000),
    .INIT_09(256'h00000000000000007FC0000000000000000000000000000000000FFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFC000000000000000000000000000000000000FF800000000000000),
    .INIT_0B(256'h0000000000000000000000003FE00000000000000000000000000000000007FF),
    .INIT_0C(256'h000003FFFFFFFFFFFF8000000000000000000000000000000000003FE0000000),
    .INIT_0D(256'hC00000000000000000000000000000000FF80000000000000000000000000000),
    .INIT_0E(256'h00000000000001FFFFFFFFFFFF0000000000000000000000000000000000007F),
    .INIT_0F(256'h000001FF8000000000000000000000000000000007FC00000000000000000000),
    .INIT_10(256'h00000000000000000000007FFFFFFFFFFC000000000000000000000000000000),
    .INIT_11(256'h00000000000003FF0000000000000000000000000000000003FF000000000000),
    .INIT_12(256'h0000000000000000000000000000003FFFFFFFFFF80000000000000000000000),
    .INIT_13(256'h000000000000000000000FFC0000000000000000000000000000000001FF8000),
    .INIT_14(256'h007FE0000000000000000000000000000000001FFFFFFFFFF000000000000000),
    .INIT_15(256'h00000000000000000000000000001FF800000000000000000000000000000000),
    .INIT_16(256'h00000000003FF0000000000000000000000000000000000FFFFFFFFFE0000000),
    .INIT_17(256'hC000000000000000000000000000000000007FE0000000000000000000000000),
    .INIT_18(256'h0000000000000000000FFC0000000000000000000000000000000007FFFFFFFF),
    .INIT_19(256'hFFFFFFFF800000000000000000000000000000000000FFC00000000000000000),
    .INIT_1A(256'h0000000000000000000000000007FE0000000000000000000000000000000003),
    .INIT_1B(256'h00000001FFFFFFFF000000000000000000000000000000000003FF0000000000),
    .INIT_1C(256'h000000000000000000000000000000000001FF80000000000000000000000000),
    .INIT_1D(256'h0000000000000000FFFFFFFE00000000000000000000000000000000000FFE00),
    .INIT_1E(256'h003FF800000000000000000000000000000000000000FFE00000000000000000),
    .INIT_1F(256'h0000000000000000000000007FFFFFFC00000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_081920_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_addra_o ,addra[14:13]}),
    .dia({open_n1690,open_n1691,open_n1692,open_n1693,open_n1694,open_n1695,open_n1696,1'b0,open_n1697}),
    .rsta(rsta),
    .doa({open_n1712,open_n1713,open_n1714,open_n1715,open_n1716,open_n1717,open_n1718,open_n1719,inst_doa_i10_000}));
  // address_offset=81920;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFC00000000000000000000000000000000FFFFFFFFFFFFFFFFFFF8FFF),
    .INIT_01(256'hFFFFBFFFFFFFFFFFFFFC00000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFF8000000000000000000000000000000007FFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000FFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000003FFFFFF),
    .INIT_05(256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000003FFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000),
    .INIT_07(256'h00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000007FFFF),
    .INIT_08(256'h001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000),
    .INIT_09(256'h0000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000),
    .INIT_0A(256'h00000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000),
    .INIT_0B(256'h000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800),
    .INIT_0C(256'hFFFFFC0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000),
    .INIT_0D(256'h000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFE000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80),
    .INIT_0F(256'hFFFFFE00000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFF800000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFC00000000000000000000000000000000000000FFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000007FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000007FFF),
    .INIT_14(256'h00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000FFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000),
    .INIT_16(256'h0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000001FFFFFFF),
    .INIT_17(256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000),
    .INIT_18(256'h0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000),
    .INIT_19(256'h000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000),
    .INIT_1A(256'h000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC),
    .INIT_1B(256'hFFFFFFFE00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000),
    .INIT_1C(256'h000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFF00000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000),
    .INIT_1E(256'hFFC00000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFF80000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_081920_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_addra_o ,addra[14:13]}),
    .dia({open_n1748,open_n1749,open_n1750,open_n1751,open_n1752,open_n1753,open_n1754,1'b0,open_n1755}),
    .rsta(rsta),
    .doa({open_n1770,open_n1771,open_n1772,open_n1773,open_n1774,open_n1775,open_n1776,open_n1777,inst_doa_i10_001}));
  // address_offset=81920;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_081920_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_addra_o ,addra[14:13]}),
    .dia({open_n1806,open_n1807,open_n1808,open_n1809,open_n1810,open_n1811,open_n1812,1'b0,open_n1813}),
    .rsta(rsta),
    .doa({open_n1828,open_n1829,open_n1830,open_n1831,open_n1832,open_n1833,open_n1834,open_n1835,inst_doa_i10_002}));
  // address_offset=90112;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000007FF0000000000000000000000000000000000000003FF800000000),
    .INIT_01(256'h000000000000000000000000000000003FFFFFF8000000000000000000000000),
    .INIT_02(256'h000000000000000001FFC0000000000000000000000000000000000000001FFC),
    .INIT_03(256'h000007FF000000000000000000000000000000001FFFFFF00000000000000000),
    .INIT_04(256'h00000000000000000000000007FF000000000000000000000000000000000000),
    .INIT_05(256'h00000000000001FFC00000000000000000000000000000001FFFFFF000000000),
    .INIT_06(256'h000000000000000000000000000000001FFC0000000000000000000000000000),
    .INIT_07(256'h00000000000000000000007FF00000000000000000000000000000000FFFFFE0),
    .INIT_08(256'h07FFFFC0000000000000000000000000000000007FF800000000000000000000),
    .INIT_09(256'h0000000000000000000000000000003FFC000000000000000000000000000000),
    .INIT_0A(256'h0000000003FFFF8000000000000000000000000000000001FFE0000000000000),
    .INIT_0B(256'h000000000000000000000000000000000000000FFF0000000000000000000000),
    .INIT_0C(256'h000000000000000001FFFF0000000000000000000000000000000007FF800000),
    .INIT_0D(256'hFE0000000000000000000000000000000000000000000003FFC0000000000000),
    .INIT_0E(256'h00000000000000000000000001FFFF000000000000000000000000000000003F),
    .INIT_0F(256'h000000FFF80000000000000000000000000000000000000000000000FFF80000),
    .INIT_10(256'h3FFE000000000000000000000000000000FFFE00000000000000000000000000),
    .INIT_11(256'h00000000000003FFE00000000000000000000000000000000000000000000000),
    .INIT_12(256'h000000000FFF8000000000000000000000000000007FFC000000000000000000),
    .INIT_13(256'h000000000000000000001FFF8000000000000000000000000000000000000000),
    .INIT_14(256'h000000000000000003FFF000000000000000000000000000003FFC0000000000),
    .INIT_15(256'h00000000000000000000000000007FFE00000000000000000000000000000000),
    .INIT_16(256'h00000000000000000000000000FFFC00000000000000000000000000003FF800),
    .INIT_17(256'h001FF8000000000000000000000000000003FFF0000000000000000000000000),
    .INIT_18(256'h00000000000000000000000000000000001FFF80000000000000000000000000),
    .INIT_19(256'h00000000000FF000000000000000000000000000001FFFC00000000000000000),
    .INIT_1A(256'h00000000000000000000000000000000000000000007FFF00000000000000000),
    .INIT_1B(256'h0000000000000000000FF000000000000000000000000000007FFF0000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000001FFFC00000000),
    .INIT_1D(256'h800000000000000000000000000FE00000000000000000000000000003FFF800),
    .INIT_1E(256'h1FFFE00000000000000000000000000000000000000000000000000000003FFF),
    .INIT_1F(256'h00000FFFF000000000000000000000000007E000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_090112_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_addra_o ,addra[14:13]}),
    .dia({open_n1864,open_n1865,open_n1866,open_n1867,open_n1868,open_n1869,open_n1870,1'b0,open_n1871}),
    .rsta(rsta),
    .doa({open_n1886,open_n1887,open_n1888,open_n1889,open_n1890,open_n1891,open_n1892,open_n1893,inst_doa_i11_000}));
  // address_offset=90112;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFF8000000000000000000000000000000000000000000007FFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000003),
    .INIT_03(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000FFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000),
    .INIT_05(256'h00000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000FFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000001F),
    .INIT_08(256'hF800003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFC00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000),
    .INIT_0B(256'h000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000),
    .INIT_0D(256'h000000000000000000000000000000000000000000000000003FFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0),
    .INIT_0F(256'hFFFFFF000000000000000000000000000000000000000000000000000007FFFF),
    .INIT_10(256'h0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF8003FFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000),
    .INIT_14(256'h000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC003FFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000),
    .INIT_16(256'h000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFC007FF),
    .INIT_17(256'hFFE007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000),
    .INIT_18(256'h000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFF00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000),
    .INIT_1A(256'h00000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFF00FFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000),
    .INIT_1C(256'h00000000000000000000000000000000000000000000000000000003FFFFFFFF),
    .INIT_1D(256'h7FFFFFFFFFFFFFFFFFFFFFFFFFF01FFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000),
    .INIT_1E(256'hE000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h000000000FFFFFFFFFFFFFFFFFFFFFFFFFF81FFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_090112_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_addra_o ,addra[14:13]}),
    .dia({open_n1922,open_n1923,open_n1924,open_n1925,open_n1926,open_n1927,open_n1928,1'b0,open_n1929}),
    .rsta(rsta),
    .doa({open_n1944,open_n1945,open_n1946,open_n1947,open_n1948,open_n1949,open_n1950,open_n1951,inst_doa_i11_001}));
  // address_offset=90112;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_090112_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_Naddra[15]_addra_o ,addra[14:13]}),
    .dia({open_n1980,open_n1981,open_n1982,open_n1983,open_n1984,open_n1985,open_n1986,1'b0,open_n1987}),
    .rsta(rsta),
    .doa({open_n2002,open_n2003,open_n2004,open_n2005,open_n2006,open_n2007,open_n2008,open_n2009,inst_doa_i11_002}));
  // address_offset=98304;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000001FFFF0000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h00000000000001FFFF00000000000000000000000003C0000000000000000000),
    .INIT_02(256'h000000000000000FFFF800000000000000000000000000000000000000000000),
    .INIT_03(256'h00000000000000000000003FFFE0000000000000000000000003C00000000000),
    .INIT_04(256'h00000000000000000000007FFFE0000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000FFFFC0000000000000000000000038000),
    .INIT_06(256'h000180000000000000000000000007FFFF000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000001FFFFC0000000000000000000),
    .INIT_08(256'h0000000000018000000000000000000000007FFFF80000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000003FFFFC0000000000),
    .INIT_0A(256'h00000000000000000000000000000000000000000007FFFF8000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000003FFFFC0),
    .INIT_0C(256'h007FFFFC0000000000000000000000000000000000000000007FFFFC00000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h00000000000FFFFFC00000000000000000000000000000000000000007FFFFE0),
    .INIT_0F(256'hFFFFFE0000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h00000000000000000000FFFFFE00000000000000000000000000000000000000),
    .INIT_11(256'h0000001FFFFFE000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h00000000000000000000000000000FFFFFF00000000000000000000000000000),
    .INIT_13(256'h00000000000007FFFFFE00000000000000000000000000000000000000000000),
    .INIT_14(256'h00000000000000000000000000000000000000FFFFFFC0000000000000000000),
    .INIT_15(256'h00000000000000000003FFFFFFE0000000000000000000000000000000000000),
    .INIT_16(256'h00000000000000000000000000000000000000000000000FFFFFFF8000000000),
    .INIT_17(256'h00000000000000000000000001FFFFFFFE000000000000000000000000000000),
    .INIT_18(256'h00000000000000000000000000000000000000000000000000000000FFFFFFFF),
    .INIT_19(256'h07FFFFFFFF0000000000000000000001FFFFFFFFC00000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h00000000003FFFFFFFFFE0000000000000000FFFFFFFFFF80000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h00000000000000000000FFFFFFFFFFFFF00000001FFFFFFFFFFFFE0000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_098304_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_addra[_o ,addra[14:13]}),
    .dia({open_n2038,open_n2039,open_n2040,open_n2041,open_n2042,open_n2043,open_n2044,1'b0,open_n2045}),
    .rsta(rsta),
    .doa({open_n2060,open_n2061,open_n2062,open_n2063,open_n2064,open_n2065,open_n2066,open_n2067,inst_doa_i12_000}));
  // address_offset=98304;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFE00000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFC3FFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000),
    .INIT_03(256'h000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFC3FFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000),
    .INIT_05(256'h000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFC7FFF),
    .INIT_06(256'hFFFE7FFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000),
    .INIT_07(256'h000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000),
    .INIT_09(256'h000000000000000000000000000000000000000000000000000003FFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000),
    .INIT_0B(256'h000000000000000000000000000000000000000000000000000000000000003F),
    .INIT_0C(256'h00000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h00000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h00000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFE000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h00000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000),
    .INIT_14(256'h000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000007FFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000FFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h000000000000000000001FFFFFFFFFFFFFFFF000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h000000000000000000000000000000000FFFFFFFE00000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_098304_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_addra[_o ,addra[14:13]}),
    .dia({open_n2096,open_n2097,open_n2098,open_n2099,open_n2100,open_n2101,open_n2102,1'b0,open_n2103}),
    .rsta(rsta),
    .doa({open_n2118,open_n2119,open_n2120,open_n2121,open_n2122,open_n2123,open_n2124,open_n2125,inst_doa_i12_001}));
  // address_offset=98304;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_098304_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_addra[_o ,addra[14:13]}),
    .dia({open_n2154,open_n2155,open_n2156,open_n2157,open_n2158,open_n2159,open_n2160,1'b0,open_n2161}),
    .rsta(rsta),
    .doa({open_n2176,open_n2177,open_n2178,open_n2179,open_n2180,open_n2181,open_n2182,open_n2183,inst_doa_i12_002}));
  // address_offset=106496;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFF80000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFF80000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h00000000000000000000000000000000000000000000000003FFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000007FFF),
    .INIT_06(256'h000000003FFFFFFFF80000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_106496_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_addra[_o ,addra[14:13]}),
    .dia({open_n2212,open_n2213,open_n2214,open_n2215,open_n2216,open_n2217,open_n2218,1'b0,open_n2219}),
    .rsta(rsta),
    .doa({open_n2234,open_n2235,open_n2236,open_n2237,open_n2238,open_n2239,open_n2240,open_n2241,inst_doa_i13_000}));
  // address_offset=106496;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_106496_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_addra[_o ,addra[14:13]}),
    .dia({open_n2270,open_n2271,open_n2272,open_n2273,open_n2274,open_n2275,open_n2276,1'b0,open_n2277}),
    .rsta(rsta),
    .doa({open_n2292,open_n2293,open_n2294,open_n2295,open_n2296,open_n2297,open_n2298,open_n2299,inst_doa_i13_001}));
  // address_offset=114688;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_114688_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_addra[_o ,addra[14:13]}),
    .dia({open_n2328,open_n2329,open_n2330,open_n2331,open_n2332,open_n2333,open_n2334,1'b0,open_n2335}),
    .rsta(rsta),
    .doa({open_n2350,open_n2351,open_n2352,open_n2353,open_n2354,open_n2355,open_n2356,open_n2357,inst_doa_i14_000}));
  // address_offset=122880;data_offset=0;depth=7680;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_130560x8_sub_122880_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({\and_addra[15]_addra[_o ,addra[14:13]}),
    .dia({open_n2386,open_n2387,open_n2388,open_n2389,open_n2390,open_n2391,open_n2392,1'b0,open_n2393}),
    .rsta(rsta),
    .doa({open_n2408,open_n2409,open_n2410,open_n2411,open_n2412,open_n2413,open_n2414,open_n2415,inst_doa_i15_000}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_1  (
    .i0(inst_doa_i2_000),
    .i1(inst_doa_i3_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_2  (
    .i0(inst_doa_i4_000),
    .i1(inst_doa_i5_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_2 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_3  (
    .i0(inst_doa_i6_000),
    .i1(inst_doa_i7_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_3 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_4  (
    .i0(inst_doa_i8_000),
    .i1(inst_doa_i9_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_4 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_5  (
    .i0(inst_doa_i10_000),
    .i1(inst_doa_i11_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_5 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_6  (
    .i0(inst_doa_i12_000),
    .i1(inst_doa_i13_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_6 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_7  (
    .i0(inst_doa_i14_000),
    .i1(inst_doa_i15_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_7 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b0/B0_0 ),
    .i1(\inst_doa_mux_b0/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b0/B0_2 ),
    .i1(\inst_doa_mux_b0/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b0/B0_4 ),
    .i1(\inst_doa_mux_b0/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_2 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b0/B0_6 ),
    .i1(\inst_doa_mux_b0/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_3 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b0/B1_0 ),
    .i1(\inst_doa_mux_b0/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b0/B1_2 ),
    .i1(\inst_doa_mux_b0/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b0/B2_0 ),
    .i1(\inst_doa_mux_b0/B2_1 ),
    .sel(addra_piped[3]),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_1  (
    .i0(inst_doa_i2_001),
    .i1(inst_doa_i3_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_2  (
    .i0(inst_doa_i4_001),
    .i1(inst_doa_i5_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_2 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_3  (
    .i0(inst_doa_i6_001),
    .i1(inst_doa_i7_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_3 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_4  (
    .i0(inst_doa_i8_001),
    .i1(inst_doa_i9_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_4 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_5  (
    .i0(inst_doa_i10_001),
    .i1(inst_doa_i11_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_5 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_6  (
    .i0(inst_doa_i12_001),
    .i1(inst_doa_i13_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_6 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_7  (
    .i0(inst_doa_i14_000),
    .i1(inst_doa_i15_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_7 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b1/B0_0 ),
    .i1(\inst_doa_mux_b1/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b1/B0_2 ),
    .i1(\inst_doa_mux_b1/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b1/B0_4 ),
    .i1(\inst_doa_mux_b1/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_2 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b1/B0_6 ),
    .i1(\inst_doa_mux_b1/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_3 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b1/B1_0 ),
    .i1(\inst_doa_mux_b1/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b1/B1_2 ),
    .i1(\inst_doa_mux_b1/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b1/B2_0 ),
    .i1(\inst_doa_mux_b1/B2_1 ),
    .sel(addra_piped[3]),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_1  (
    .i0(inst_doa_i2_002),
    .i1(inst_doa_i3_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_2  (
    .i0(inst_doa_i4_002),
    .i1(inst_doa_i5_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_2 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_3  (
    .i0(inst_doa_i6_002),
    .i1(inst_doa_i7_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_3 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_4  (
    .i0(inst_doa_i8_002),
    .i1(inst_doa_i9_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_4 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_5  (
    .i0(inst_doa_i10_002),
    .i1(inst_doa_i11_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_5 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_6  (
    .i0(inst_doa_i12_002),
    .i1(inst_doa_i13_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_6 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_7  (
    .i0(inst_doa_i14_000),
    .i1(inst_doa_i15_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_7 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b2/B0_0 ),
    .i1(\inst_doa_mux_b2/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b2/B0_2 ),
    .i1(\inst_doa_mux_b2/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b2/B0_4 ),
    .i1(\inst_doa_mux_b2/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_2 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b2/B0_6 ),
    .i1(\inst_doa_mux_b2/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_3 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b2/B1_0 ),
    .i1(\inst_doa_mux_b2/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b2/B1_2 ),
    .i1(\inst_doa_mux_b2/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b2/B2_0 ),
    .i1(\inst_doa_mux_b2/B2_1 ),
    .sel(addra_piped[3]),
    .o(doa[2]));

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

